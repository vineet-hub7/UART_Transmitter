`timescale 1ns / 1ps

module baud_gen_test(

    );
endmodule
